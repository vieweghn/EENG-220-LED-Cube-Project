//module LED_Matrix():

	