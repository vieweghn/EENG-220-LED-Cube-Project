module snpnoinoinpom
